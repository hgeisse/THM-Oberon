//
// risc5cpu.v -- the RISC5 CPU
//


`timescale 1ns/1ps
`default_nettype none


module risc5cpu(
    input clk,
    input rst);

endmodule
