//
// risc5top.v -- RISC5 toplevel description
//


`timescale 1ns/1ps
`default_nettype none


module risc5top(
    input clk_in,
    input rst_in_n);

endmodule
