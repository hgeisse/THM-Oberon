//
// PS2Dev.v -- PS/2 Interface
//


`timescale 1ns / 1ps
`default_nettype none


module PS2Dev();

endmodule
