//
// cpu.v -- RISC5 CPU
//


`timescale 1ns / 1ps
`default_nettype none


module cpu(clk, rst);
    input clk;
    input rst;

  //
  // IF stage
  //

  //
  // ID stage
  //

  //
  // EX stage
  //

  //
  // MEM stage
  //

  //
  // WB stage
  //

endmodule
