//
// RS232Dev.v -- Serial line
//


`timescale 1ns / 1ps
`default_nettype none


module RS232Dev();

endmodule
